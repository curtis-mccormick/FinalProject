module outfunction #(
    parameters
) (
    //seed
    //initial seed: 0412_6424_0034_3C28
    //next seed:    0006_7E60_3824_042C
    //seed
    assign grid = 64'h0412_6424_0034_3C28;


    datapath(grid, grid_evolve );

    grid_evolve [7:0] 

);
    
endmodule